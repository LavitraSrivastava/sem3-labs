`timescale 1ns/1ns
`include "Encoder16_4.v"

module Encoder16_4_tb;
    reg [15:0] w;
    wire [3:0] y;
    wire z;


Encoder16_4 q(w, y, z);

initial begin
        $dumpfile("Encoder16_4_tb.vcd");
        $dumpvars(0, Encoder16_4_tb);


        w = 16'b0000000000000000; #20;
        w = 16'b0000000000000010; #20;
        w = 16'b0000000000000100; #20;
        w = 16'b0000000000001000; #20;
        w = 16'b0000000000010000; #20;
        w = 16'b0000000000100000; #20;
        w = 16'b0000000001000000; #20;
        w = 16'b0000000010000000; #20;
        w = 16'b0000000100000000; #20;
        w = 16'b0000001000000000; #20;
        w = 16'b0000010000000000; #20;
        w = 16'b0000100000000000; #20;
        w = 16'b0001000000000000; #20;
        w = 16'b0010000000000000; #20;
        w = 16'b0100000000000000; #20;
        w = 16'b1000000000000000; #20;

        $display("Test Complete");
    end
endmodule
