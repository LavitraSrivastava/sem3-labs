`timescale 1ns/1ns
`include "PEn16to4.v"

module PEn16to4_tb();
reg [15:0]w;
wire [3:0]y;
wire z;

PEn16to4 p2(w,y,z);
initial begin
$dumpfile("PEn16to4_tb.vcd");
$dumpvars(0, PEn16to4_tb);

w=16'b1000000000000000;#20;
w=16'b0100000000000000;#20;
w=16'b0010000000000000;#20;
w=16'b0001000000000000;#20;
w=16'b0000100000000000;#20;
w=16'b0000010000000000;#20;
w=16'b0000001000000000;#20;
w=16'b0000000100000000;#20;
w=16'b0000000010000000;#20;
w=16'b0000000001000000;#20;
w=16'b0000000000100000;#20;
w=16'b0000000000010000;#20;
w=16'b0000000000001000;#20;
w=16'b0000000000000100;#20;
w=16'b0000000000000010;#20;
w=16'b0000000000000001;#20;
w=16'b0000000000000000;#20;

$display("Test complete");
end
endmodule
