module FA_dec2to4(en,w,y);
input en;
input [1
